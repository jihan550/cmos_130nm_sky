** sch_path: /home/jihan/projects/buffer/untitled.sch
**.subckt untitled
XM1 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM2 Vout Vin GND VDD sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
Vdd VDD GND 1.8
Vin Vin GND 0
**** begin user architecture code

.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.option wnflag=1


.dc Vin 0 1.8 0.01
.save all

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
